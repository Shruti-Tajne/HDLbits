// Question 2. Zero - https://hdlbits.01xz.net/wiki/Zero

module top_module ( output zero );
	
	assign zero = 1'b0;
	
endmodule

//Watch video for explanation: https://www.youtube.com/watch?v=4ynX6o0Zznw
