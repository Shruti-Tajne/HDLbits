//Question 3.Wire - https://hdlbits.01xz.net/wiki/Wire

module top_module( input in, output out );
	
	assign out = in;
	// Note that wires are directional, so "assign in = out" is not equivalent.
	
endmodule

