// Question 6. Andgate - https://hdlbits.01xz.net/wiki/Andgate

module top_module( 
    input a, 
    input b, 
    output out );
    
    assign out = a&b;

endmodule
